`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/12/2018 10:42:11 AM
// Design Name: 
// Module Name: counter_ip
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

(* use_dsp48 = "no" *)
module counter_ip(
    input clk,
    input enable,
    input up_dn,
    input reset,
    output reg [7:0] count
    );
    
    
    
endmodule
