

module comparator_dataflow(v,z);
input [3:0]v;
output z; 

assign = v[ ] 
endmodule
